module dummy_sender();

endmodule
