module dummy_receiver();



endmodule
